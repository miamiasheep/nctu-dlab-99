`timescale 1ns / 1ps
module word(
	output word,
	input [3:0] row, col,
	input [1:0] select
);
reg [15:0] line[15:0];

integer i;
always @(*)
begin
	if (select == 1) begin
		line[0] = 16'b0000000000000000;
		line[1] = 16'b0000000000000000;
		line[2] = 16'b0000111111110000;
		line[3] = 16'b0001111111111000;
		line[4] = 16'b0011100000011100;
		line[5] = 16'b0111000000001110;
		line[6] = 16'b0111000000001110;
		line[7] = 16'b0111000000001110;
		line[8] = 16'b0111000000001110;
		line[9] = 16'b0111000000001110;
		line[10] =16'b0111000000001110;
		line[11] =16'b0111000000001110;
		line[12] =16'b0111000000001110;
		line[13] =16'b0011111111111100;
		line[14] =16'b0001111111111000;
		line[15] =16'b0000000000000000;
	end else if (select == 2) begin
		line[0] = 16'b0000000000000000;
		line[1] = 16'b1110000000000111;
		line[2] = 16'b0111000000001110;
		line[3] = 16'b0011100000011100;
		line[4] = 16'b0001110000111000;
		line[5] = 16'b0000111001110000;
		line[6] = 16'b0000011111100000;
		line[7] = 16'b0000001111000000;
		line[8] = 16'b0000001111000000;
		line[9] = 16'b0000011111100000;
		line[10] =16'b0000111001110000;
		line[11] =16'b0001110000111000;
		line[12] =16'b0011100000011100;
		line[13] =16'b0111000000001110;
		line[14] =16'b1110000000000111;
		line[15] =16'b0000000000000000;
	end else for (i=0; i<16; i=i+1)
		line[i] = 16'b0;
end

assign word = (select == 0) ? 1'b0 : (line[row] >> (~col)) % 2;

endmodule
